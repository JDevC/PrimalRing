�}q (X   Coinsq]q(KKdeX   Energyq]q(KdKdeX   Lifeq]q(KRKdeX   Levelq}q(X   IDq	X   The RINGq
X	   PositionYqM�X	   PositionXqMuX   NameqX   Playerqu.